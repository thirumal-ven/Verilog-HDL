module gates_tb;
reg a,b;
wire c,d,e,f;

gates u1 


























































++














































































































































































































































































































































































































































































































































































a,b,c,d,e,f);

initial
begin
a=0;b=0;
#10 a=1'b0;b=1'b0;
#10 a=1'b0;b=1'b1;
#10 a=1'b1;b=1'b0;
#10 a=1'b1;b=1'b1;
#10 $finish;

end
endmodule
+