module mux81_tb ;
reg [7:0]i;
reg [2:0]s;
wire y;
mux81 u1 (i,s,y);
initial
begin
#10 s[0]=1'b0;s[1]=1'b0;s[2]=1'b0;
#10 s[0]=1'b0;s[1]=0;s[2]=1'b0;i[0]=1'b1;i[0]=1'b0;i[2]=1'b0;i[3]=1'b0;i[4]=1'b0;i[5]=1'b0;i[6]=1'b0;i[7]=1'b0;
#10 s[0]=1'b0;s[1]=0;s[2]=1'b1;i[1]=1'b1;i[2]=1'b0;i[0]=1'b0;i[3]=1'b0;i[4]=1'b0;i[5]=1'b0;i[6]=1'b0;i[7]=1'b0;
#10 s[0]=1'b0;s[1]=1;s[2]=1'b0;i[2]=1'b1;i[1]=1'b0;i[3]=1'b0;i[0]=1'b0;i[4]=1'b0;i[5]=1'b0;i[6]=1'b0;i[7]=1'b0;
#10 s[0]=1'b0;s[1]=1;s[2]=1'b1;i[3]=1'b1;i[1]=1'b0;i[2]=1'b0;i[4]=1'b0;i[0]=1'b0;i[5]=1'b0;i[6]=1'b0;i[7]=1'b0;
#10 s[0]=1'b1;s[1]=0;s[2]=1'b0;i[4]=1'b1;i[1]=1'b0;i[2]=1'b0;i[3]=1'b0;i[5]=1'b0;i[0]=1'b0;i[6]=1'b0;i[7]=1'b0;
#10 s[0]=1'b1;s[1]=0;s[2]=1'b1;i[5]=1'b1;i[1]=1'b0;i[2]=1'b0;i[3]=1'b0;i[4]=1'b0;i[6]=1'b0;i[0]=1'b0;i[7]=1'b0;
#10 s[0]=1'b1;s[1]=1;s[2]=1'b0;i[6]=1'b1;i[1]=1'b0;i[2]=1'b0;i[3]=1'b0;i[4]=1'b0;i[5]=1'b0;i[7]=1'b0;i[0]=1'b0;
#10 s[0]=1'b1;s[1]=1;s[2]=1'b1;i[7]=1'b1;i[1]=1'b0;i[2]=1'b0;i[3]=1'b0;i[4]=1'b0;i[5]=1'b0;i[6]=1'b0;i[0]=1'b0;
#10 $finish ;
end 
endmodule
